../lib/python3.12
../lib/python3.12/lib-dynload
../lib/python3.12/site-packages 
../lib/python3.12/dist-packages 
../lib/python312.zip 
